package i2c_enum;
typedef enum bit {wr,rd}i2c_op_t ;
endpackage