
typedef enum bit {wr,rd}i2c_op_t ; 

