b0VIM 7.4      ��9b&1�
�(  smamidi                                 grendel29.ece.ncsu.edu                  ~smamidi/ECE745/ece745_projects/project_benches/proj_1/testbench/top.sv                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                     ���������       �                             K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     �       �  �  �  �  �  �  �  a  @          �  �  �  �  �  �  w  m  N  /      �  �  �  |  i  h  `  P  F  5  1  0  �  �  �  �  �  �  �  �  P        �  �  �  �  h            �
  �
  �
  �
  g
  N
  M
  @
  4
  3
  2
   
  
  �	  �	  �	  �	  {	  k	  g	  B	  	  �  �  �  �  �  �  k  F  @  0  ,    �  �  �  �  �  �  o  I  C  3  /  
    �  �  �  �  �  x  w  v  u  n  m  E    �  �  �  �  �  �  h  B  <  ,  (    �  �  �  �  ~  z  U  C  =    �  �  �  �  �  �  Y  U  -      �  �  �  �  �                     wb_bus.master_read(2'h01,receiving_data); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7])|| (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx011); end $display("Read Data is : %d",receiving_data); wb_bus.master_read(2'h01,receiving_data); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7])|| (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx010); begin for(i=0;i<31;i++) wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7])|| (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx001); wb_bus.master_write(2'h01,8'h45); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx100); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx110); wb_bus.master_write(2'h01,8'b00000101); wb_bus.master_write(2'h00,8'b11xxxxxx);  //READ    wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin  while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx101); end wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx001); wb_bus.master_write(2'h01,i); for(int i=0; i<32; i++) begin end @(posedge clk); begin while(!(wb_bus.dat_o[6])) wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7])|| (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx001); wb_bus.master_write(2'h01,8'h44); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx100); wb_bus.master_read(2'h02,cmdr_data); end @(posedge clk); begin while(!(wb_bus.dat_o[7]) || (!(irq))) wb_bus.master_write(2'h02,8'bxxxxx110); wb_bus.master_write(2'h01,8'b00000101); wb_bus.master_write(2'h00,8'b11xxxxxx);  //WRITE execution   write_i=64; int write_i;  bit[7:0] receiving_data; reg [WB_DATA_WIDTH-1:0]cmdr_data;  initial begin :test_flow // Define the flow of the simulation // ****************************************************************************    end   //$display("addr=%0xh, data=%0xh, Write enable = %d",adr,dat_wr_o,we);   wb_bus.master_monitor(.addr(addrwr),.data(datwr),.we(wen));  bit wen;  bit [WB_ADDR_WIDTH-1:0] addrwr;  bit [WB_DATA_WIDTH-1:0] datwr; begin: wb_monitoring initial   // Monitor Wishbone bus and display transfers in the transcript // ****************************************************************************  end #113 rst=1'b0; begin : rst_gen initial  // Reset generator // ****************************************************************************  end     #5 clk=~clk;   forever begin : clk_gen initial  // Clock generator // **************************************************************************** int temp1=0; i2c_op_t op_top; bit [7:0]i2c_read_data[]; int i; bit [WB_ADDR_WIDTH-1:0] data_out[]; tri  [NUM_I2C_BUSSES-1:0] sda; tri  [NUM_I2C_BUSSES-1:0] scl; wire irq; wire [WB_DATA_WIDTH-1:0] dat_rd_i; wire [WB_DATA_WIDTH-1:0] dat_wr_o; wire [WB_ADDR_WIDTH-1:0] adr; tri1 ack; wire we; wire stb; wire cyc; bit  rst = 1'b1; bit  clk;  parameter int NUM_I2C_BUSSES = 1; parameter int WB_DATA_WIDTH = 8; parameter int i2c_DATA_WIDTH = 8; parameter int WB_ADDR_WIDTH = 2; parameter int i2c_ADDR_WIDTH = 7; module top();   import i2c_pkg ::*; `timescale 1ns / 10ps ad  �  ,	             �  �  �  |  +  �  �  E  �  �  $  �  v    �  �  �  M  !  �
  �
  
  $
  �	  k	  ?	  :	  9	  8	  .	  -	  ,	  +	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    endmodule     );     // ------------------------------------     .sda_o(sda)          //   out std_logic_vector(0 to g_bus_num - 1)  -- I2C Data outputs     .scl_o(scl),         //   out std_logic_vector(0 to g_bus_num - 1); -- I2C Clock outputs     .sda_i(sda),         // in    std_logic_vector(0 to g_bus_num - 1); -- I2C Data inputs     .scl_i(scl),         // in    std_logic_vector(0 to g_bus_num - 1); -- I2C Clock inputs     // -- I2C interfaces:     // ------------------------------------     // ------------------------------------     .irq(irq),           //   out std_logic;                            -- Interrupt request     // -- Interrupt request:     // ------------------------------------     // ------------------------------------     .dat_o(dat_rd_i),    //   out std_logic_vector(7 downto 0);         -- Data output     .dat_i(dat_wr_o),    // in    std_logic_vector(7 downto 0);         -- Data input     .we_i(we),           // in    std_logic;                            -- Write enable     .adr_i(adr),         // in    std_logic_vector(1 downto 0);         -- Low bits of Wishbone address     .ack_o(ack),         //   out std_logic;                            -- Acknowledge output     .stb_i(stb),         // in    std_logic;                            -- Slave selection     .cyc_i(cyc),         // in    std_logic;                            -- Valid bus cycle indication     // -------------     .rst_i(rst),         // in    std_logic;                            -- Synchronous reset (active high)     .clk_i(clk),         // in    std_logic;                            -- Clock     // -- Wishbone signals:     // ------------------------------------   ( \work.iicmb_m_wb(str) #(.g_bus_num(NUM_I2C_BUSSES)) DUT 